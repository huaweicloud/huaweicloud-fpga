//
//------------------------------------------------------------------------------
//     Copyright (c) 2017 Huawei Technologies Co., Ltd. All Rights Reserved.
//
//     This program is free software; you can redistribute it and/or modify
//     it under the terms of the Huawei Software License (the "License").
//     A copy of the License is located in the "LICENSE" file accompanying 
//     this file.
//
//     This program is distributed in the hope that it will be useful,
//     but WITHOUT ANY WARRANTY; without even the implied warranty of
//     MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the
//     Huawei Software License for more details. 
//------------------------------------------------------------------------------


`ifndef _TB_PKG_SVH_
`define _TB_PKG_SVH_

// package tb_pkg;

// ./test/tb_env.sv
`include "tb_env.sv"
// ./test/tb_test.sv
`include "tb_test.sv"

// endpackage

// ./tb_top.sv
// `include "tb_top.sv"

`endif // _TB_PKG_SVH_

